import uvm_pkg::*;

module tb_top();
  initial begin
    run_test();
  end
endmodule
