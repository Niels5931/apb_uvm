
package pk_apb;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "apb_common.svh"
  `include "cl_apb_seq_item.svh"

endpackage : pk_apb
