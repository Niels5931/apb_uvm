interface if_clk#(
  parameter NUM_OF_CLOCKS = 1
) (
  input logic PCLK,
  input logic PRESETn
);

endinterface : if_clk

