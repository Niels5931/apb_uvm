package pk_apb_vseqs;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "cl_apb_tb_simple_vseq.svh"

endpackage : pk_apb_vseqs
