package pk_apb_tb;

  `include "cl_uvm_simple_test.svh"

endpackage : pk_apb_tb
