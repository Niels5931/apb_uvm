package pk_apb_test;

  `include "uvm_macros.svh"
  `include "cl_apb_tb_simple_test.svh"

endpackage : pk_apb_test
