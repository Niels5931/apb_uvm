typedef enum{
  RD = 1'b0,
  WR = 1'b1
} op_type;
