
package pk_apb;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "apb_common.svh"
  `include "cl_apb_seq_item.svh"
  `include "cl_apb_seq_lib.svh"
  `include "cl_apb_config.svh"
  `include "cl_apb_driver_base.svh"
  `include "cl_apb_driver_manager.svh"
  `include "cl_apb_agent.svh"

endpackage : pk_apb
