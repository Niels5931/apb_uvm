package pk_apb_tests;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "cl_apb_tb_simple_test.svh"
  `include "cl_uvm_simple_test.svh"

endpackage : pk_apb_tests
