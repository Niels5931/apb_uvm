package pk_apb_tb;
  import uvm_pkg::*;
  import pk_apb::*;
  `include "uvm_macros.svh"
  `include "cl_apb_tb_vseqr.svh"
  `include "cl_apb_tb_config.svh"
  `include "cl_apb_tb_env.svh"
  `include "cl_apb_tb_base_vseq.svh"
  `include "cl_apb_tb_base_test.svh"

endpackage : pk_apb_tb
