import pkg_uvm::*;

package pk_apb_tb;

  `include "uvm_macros.svh"
  `include "cl_apb_tb_vseqr.svh"
  `include "cl_apb_tb_env.svh"

endpackage : pk_apb_tb
